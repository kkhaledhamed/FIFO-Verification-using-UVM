package FIFO_shared_pkg;

	// Counters to be used in scoreboard
	integer correct_count = 0;
	integer error_count = 0;

endpackage 